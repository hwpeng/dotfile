module  
(
	input clk_i
	,input rst_i

);

endmodule
